--Instruction Register Block