--Memory Interface Block