-- Operational decode block for Control Unit