--Arithmetic Logic Unit Block