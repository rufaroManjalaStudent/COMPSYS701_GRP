-- sys_clock.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sys_clock is
	port (
		clk : out std_logic   -- clk.clk
	);
end entity sys_clock;

architecture rtl of sys_clock is
	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

begin

	clock_source_0 : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50,
			CLOCK_UNIT => 1000000
		)
		port map (
			clk => clk  -- clk.clk
		);

end architecture rtl; -- of sys_clock
