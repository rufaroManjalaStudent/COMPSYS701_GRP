library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity resetGen is
	port (
	);
end entity resetGen;

architecture behaviour of resetGen is
begin

end architecture behaviour;