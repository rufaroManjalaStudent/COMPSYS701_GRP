
module sys_clock (
	clk);	

	output		clk;
endmodule
