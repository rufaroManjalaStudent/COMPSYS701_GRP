--Control Unit sub-top-level design
