-- Operational decode block for Control Unit
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OpDec is
    port(
        state       : in std_logic_vector(2 downto 0);
    )

end entity;

architecture behaviour of OpDec is
    --signal declaration
    begin 

end architecture;